module alu #(parameter WIDTH = 32) (
    input       [WIDTH-1:0] a, b,       // operands
    input       [2:0] alu_ctrl,         // ALU control
    input       funct7b5, funct3,       // funct7[5] and funct3[0]
    output reg  [WIDTH-1:0] alu_out,    // ALU output
    output      Zero                    // zero flag
);

always @(*) begin
    case (alu_ctrl)
        3'b000:  alu_out <= a + b;           // ADD/ADDI
        3'b001:  alu_out <= a - b;           // SUB/SUBI
        3'b010:  alu_out <= $signed(a) < $signed(b) ? 1 : 0; // SLT (signed comparison)
        3'b110:  alu_out <= a < b ? 1 : 0;   // SLTU (unsigned comparison)
        3'b100:  alu_out <= a ^ b;           // XOR/XORI
        3'b101: begin                        // Shift operations
            if (funct7b5) alu_out <= $signed(a) >>> b[4:0];   // SRA/SRAI (arithmetic shift)
            else alu_out <= a >> b[4:0];                      // SRL/SRLI (logical shift)
        end
        3'b011:  alu_out <= a | b;           // OR/ORI
        3'b111:  alu_out <= a << b[4:0];     // SLL/SLLI (Shift Left Logical)
        default: alu_out <= 0;               // Default case (no operation)
    endcase
end

assign Zero = (alu_out == 0) ? 1'b1 : 1'b0;               // Zero flag

endmodule

